
module lab1 (
	clk_clk,
	led_export,
	reset_reset_n,
	bouton_export);	

	input		clk_clk;
	output	[7:0]	led_export;
	input		reset_reset_n;
	input	[7:0]	bouton_export;
endmodule
